module pcie_ltssm_sm (
  input  logic clk,
  input  logic reset,
  output logic link_up
);

endmodule
