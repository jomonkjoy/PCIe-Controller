module byte_striping #(
) (
);

endmodule

module byte_striping #(
) (
);

endmodule
